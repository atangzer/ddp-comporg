`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:22:30 03/14/2020 
// Design Name: 
// Module Name:    Counter_x 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Counter_x(input clk,			//io_clk			    input rst,			    input clk0,			//clk_div[7],??U8			    input clk1,			// clk_div[10],??U8			    input clk2,			//clk_div[10],??U8			    input counter_we,		//??????,??U4			    input [31:0] counter_val,        //???????,??U4			    input [1:0] counter_ch,	           //???????,??U7								    output counter0_OUT,		//???U4			    output counter1_OUT,		 //???U4			    output counter2_OUT,		 //???U4			    output [31:0] counter_out	 //???U4			   );endmodule


endmodule
